module top_module(
    input a,b,
    output y
);
    assign y = a & b;
endmodule
