module and2_prim (
    input  a,
    input  b,
    output y
);
    // TODO: instantiate the built-in AND gate primitive
    // and <instance_name> ( <out>, <in1>, <in2> );
    and a1(y,a,b);
endmodule
