module selector3(
    input [7:0]a,b,c,
    input [1:0]sel,
    output reg [7:0]y
);

always@(*)begin
    if(sel==2'b00)
        y = a;
    else if(sel==2'b01)
        y = b;
    else if(sel==2'b10)
        y = c;
    else
        y = 8'h00;
end
endmodule
