module top_module(
    input a,
    output y
);
    assign y = ~a;
endmodule
