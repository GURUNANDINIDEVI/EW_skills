// Connect one input a to three outputs y1, y2, and y3 using wires. All outputs must always match the input.

// Requirements:

// Module Name: top_module
// Inputs: a (1-bit)
// Outputs: y1, y2, y3 (1-bit each)
module top_module(
    input a,
    output y1,y2,y3
);
    assign y1 = a;
    assign y2 = a;
    assign y3 = a;

endmodule
